`timescale 1ns / 1ps

/*******************************************************************
*
* Module: shifter0.v
* Project: femtorv32
* Authors: Mahinour Abdelgawad mahinourabdelgawad@aucegypt.edu
           Joudy ElGayar Joudyelgayar@aucegypt.edu
           
* Description:
*
* Change history: 7/11/2025 - Created module 
* 
*
**********************************************************************/

module shifter0(

    );
endmodule

