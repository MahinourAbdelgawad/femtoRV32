`timescale 1ns / 1ps

module InstMem (input [5:0] addr, output [31:0] data_out);
reg [31:0] mem [0:63];

initial begin : init_rom
integer i;
for (i = 0; i < 64; i = i + 1) mem[i] = 32'h00000013; // (ADDI x0,x0,0)
mem[0] = 32'h00000093; // ADDI x1,x0,0
mem[1] = 32'h00108113; // ADDI x2,x1,1
mem[2] = 32'h00210193; // ADDI x3,x2,2
mem[3] = 32'h00318213; // ADDI x4,x3,3
mem[10]= 32'h00b50633; // ADD x12,x10,x11 
end

    initial begin
    
    //Exp 1
//        mem[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
//        mem[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
//        mem[2]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
//        mem[3]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
//        mem[4]=32'b0_000000_00011_00100_000_0100_0_1100011; //beq x4, x3, 4
//        mem[5]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2 skip
//        mem[6]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
//        mem[7]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
//        mem[8]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
//        mem[9]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
//        mem[10]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
//        mem[11]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
//        mem[12]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1


        // Exp 2
//        mem[0] = 32'b00000000000000000010000010000011; // lw x1, 0(x0)
//        mem[1] = 32'b00000000010000000010000100000011; // lw x2, 4(x0)
//        mem[2] = 32'b00000000100000000010000110000011; // lw x3, 8(x0)
//        mem[3] = 32'b00000000000100010000000100110011; // add x2, x2, x1
//        mem[4] = 32'b01000000001100001000000010110011; // sub x1, x1, x3
//        mem[5] = 32'b00000000000000001000000101100011; // beq x1, x0, exit
//        mem[6] = 32'b11111110000000000000110111100011; // beq x0, x0, loop
//        mem[7] = 32'b00000000001000000010011000100011; // sw x2, 12(x0)


        // B-Type Testing
        mem[0]  = 32'h00500093; // ADDI x1, x0, 5
        mem[1]  = 32'h00500113; // ADDI x2, x0, 5
        mem[2]  = 32'h00300193; // ADDI x3, x0, 3
        mem[3]  = 32'h00208663; // BEQ x1, x2, +8
        mem[4]  = 32'h00309663; // BNE x1, x3, +8
        mem[5]  = 32'h0011C663; // BLT x3, x1, +8
        mem[6]  = 32'h0011D663; // BGE x3, x1, +8
        mem[7]  = 32'h0011E663; // BLTU x3, x1, +8
        mem[8]  = 32'h0011F663; // BGEU x3, x1, +8
        mem[9]  = 32'h00900213; // ADDI x4, x0, 9

 
    end 
    
    
assign data_out = mem[addr];
endmodule
