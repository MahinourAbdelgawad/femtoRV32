`timescale 1ns / 1ps

module InstMem (input [5:0] addr, output [31:0] data_out);
reg [31:0] mem [0:63];


//initial begin : init_rom
//  integer i;
//  for (i = 0; i < 64; i = i + 1) mem[i] = 32'h00000013; // NOP (ADDI x0,x0,0)

//  // Load values from Data Memory
//  mem[0]  = 32'b000000000000_00000_010_00001_0000011; // lw x1, 0(x0)  -> 5
//  mem[1]  = 32'b000000000100_00000_010_00010_0000011; // lw x2, 4(x0)  -> 5
//  mem[2]  = 32'b000000001000_00000_010_00011_0000011; // lw x3, 8(x0)  -> 3
//  mem[3]  = 32'b000000001100_00000_010_00100_0000011; // lw x4, 12(x0) -> 9

//  // --- BEQ Test ---
//  mem[4]  = 32'b0000000_00010_00001_000_01000_1100011; // beq x1, x2, +8  (should take)
//  mem[5]  = 32'b0000000_00011_00001_000_00000_0110011; // add x0, x1, x3  (skipped)
//  mem[6]  = 32'b0000000_00010_00001_000_00101_0110011; // add x5, x1, x2  (target)

//  // --- BNE Test ---
//  mem[7]  = 32'b0000000_00011_00001_001_01000_1100011; // bne x1, x3, +8  (should take)
//  mem[8]  = 32'b0000000_00001_00001_000_00110_0110011; // add x6, x1, x1  (skipped)
//  mem[9]  = 32'b0000000_00101_00001_000_00111_0110011; // add x7, x1, x5  (target)

//  // --- BLT Test ---
//  mem[10] = 32'b0000000_00001_00011_100_01000_1100011; // blt x3, x1, +8  (true, 3<5)
//  mem[11] = 32'b0000000_00011_00001_000_01000_0110011; // add x8, x1, x3  (skipped)
//  mem[12] = 32'b0000000_00011_00001_000_01001_0110011; // add x9, x1, x3  (target)

//  // --- BGE Test ---
//  mem[13] = 32'b0000000_00011_00001_101_01000_1100011; // bge x3, x1, +8  (false, 3>=5 false)
//  mem[14] = 32'b0000000_00011_00001_000_01010_0110011; // add x10, x1, x3 (executed)
//  mem[15] = 32'b0000000_00011_00001_000_01011_0110011; // add x11, x1, x3 (skipped if branch taken)

//  // --- BLTU Test (unsigned less than) ---
//  mem[16] = 32'b0000000_00001_00011_110_01000_1100011; // bltu x3, x1, +8 (true, 3<5 unsigned)
//  mem[17] = 32'b0000000_00011_00001_000_01100_0110011; // add x12, x1, x3 (skipped)
//  mem[18] = 32'b0000000_00011_00001_000_01101_0110011; // add x13, x1, x3 (target)

//  // --- BGEU Test (unsigned greater or equal) ---
//  mem[19] = 32'b0000000_00001_00011_111_01000_1100011; // bgeu x3, x1, +8 (false)
//  mem[20] = 32'b0000000_00011_00001_000_01110_0110011; // add x14, x1, x3 (executed)
//  mem[21] = 32'b0000000_00011_00001_000_01111_0110011; // add x15, x1, x3 (skipped if taken)
//end


initial begin : init_rom
integer i;
for (i = 0; i < 64; i = i + 1) mem[i] = 32'h00000013; // (ADDI x0,x0,0)
mem[0] = 32'h00000093; // ADDI x1,x0,0
mem[1] = 32'h00108113; // ADDI x2,x1,1
mem[2] = 32'h00210193; // ADDI x3,x2,2
mem[3] = 32'h00318213; // ADDI x4,x3,3
mem[10]= 32'h00b50633; // ADD x12,x10,x11 
end

    initial begin
    
//          mem[0]=32'b111111111011_00000_000_00001_0010011; 
//    //Exp 1
//        mem[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
//        mem[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
//        mem[2]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
//        mem[3]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
//        mem[4]=32'b0_000000_00011_00100_000_0100_0_1100011; //beq x4, x3, 4
//        mem[5]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2 skip
//        mem[6]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
//        mem[7]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
//        mem[8]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
//        mem[9]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
//        mem[10]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
//        mem[11]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
//        mem[12]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1



        // Exp 2
//        mem[0] = 32'b00000000000000000010000010000011; // lw x1, 0(x0)
//        mem[1] = 32'b00000000010000000010000100000011; // lw x2, 4(x0)
//        mem[2] = 32'b00000000100000000010000110000011; // lw x3, 8(x0)
//        mem[3] = 32'b00000000000100010000000100110011; // add x2, x2, x1
//        mem[4] = 32'b01000000001100001000000010110011; // sub x1, x1, x3
//        mem[5] = 32'b00000000000000001000000101100011; // beq x1, x0, exit
//        mem[6] = 32'b11111110000000000000110111100011; // beq x0, x0, loop
//        mem[7] = 32'b00000000001000000010011000100011; // sw x2, 12(x0)


//        // B-Type Testing
//        mem[0]  = 32'h00500093; // ADDI x1, x0, 5
//        mem[1]  = 32'h00500113; // ADDI x2, x0, 5
//        mem[2]  = 32'h00300193; // ADDI x3, x0, 3
//        mem[3]  = 32'h00208463; // BEQ  x1, x2, +8
//        mem[4]  = 32'h00309463; // BNE  x1, x3, +8
//        mem[5]  = 32'h0011C463; // BLT  x3, x1, +8
//        mem[6]  = 32'h0011D463; // BGE  x3, x1, +8
//        mem[7]  = 32'h0011E463; // BLTU x3, x1, +8
//        mem[8]  = 32'h0011F463; // BGEU x3, x1, +8
//        mem[9]  = 32'h00900213; // ADDI x4, x0, 9

    // J Type Testing
//    mem[0]  = 32'h00000013; // NOP (ADDI x0, x0, 0)
//    mem[1]  = 32'h004000EF; // JAL  x1, +4  --> jump to mem[3], x1 = PC+4 = 8
//    mem[2]  = 32'h00000013; // NOP (should be skipped)
//    mem[3]  = 32'h00800113; // ADDI x2, x0, 8
//    mem[4]  = 32'h00008167; // JALR x3, x1, 0  --> jump to x1 (return address from first JAL)
//    mem[5]  = 32'h00000013; // NOP (should be skipped if JALR works)
//    mem[6]  = 32'h00A00293; // ADDI x5, x0, 10 (check sequential execution after jump)
//    mem[7]  = 32'h00000013; // NOP

    // I Type Testing
//    mem[0] = 32'h00500093; // ADDI x1, x0, 5       ; x1 = 5
//    mem[1] = 32'h00308113; // ADDI x2, x1, 3       ; x2 = x1 + 3 = 8
//    mem[2] = 32'h00210213; // SLTI x4, x2, 2       ; x4 = (x2<2)?1:0 = 0
//    mem[3] = 32'h00211213; // SLTIU x4, x2, 2      ; x4 = (x2<2)?1:0 unsigned = 0
//    mem[4] = 32'h00312413; // XORI x8, x2, 3       ; x8 = x2 ^ 3 = 8 ^ 3 = 11
//    mem[5] = 32'h00113613; // ORI x12, x2, 1       ; x12 = x2 | 1 = 9
//    mem[6] = 32'h00114613; // ANDI x12, x2, 1      ; x12 = x2 & 1 = 0
//    mem[7] = 32'h00115513; // SLLI x10, x2, 1      ; x10 = x2 << 1 = 16
//    mem[8] = 32'h00116513; // SRLI x10, x2, 1      ; x10 = x2 >> 1 = 4
//    mem[9] = 32'h40117513; // SRAI x10, x2, 1      ; x10 = arithmetic right shift x2 >> 1 = 4
//    mem[10]= 32'h00008067; // JALR x1, x0, 0       ; PC = x0 + 0 = 0, test JALR

        mem[0] = 32'h00500093; // ADDI  x1, x0, 5       ; x1 = 5
        mem[1] = 32'h00308113; // ADDI  x2, x1, 3       ; x2 = x1 + 3 = 8
        mem[2] = 32'h00210213; // SLTI  x4, x2, 2       ; x4 = (x2<2)?1:0 = 0
        mem[3] = 32'h00211213; // SLTIU x4, x2, 2       ; x4 = (x2<2)?1:0 unsigned = 0
        mem[4] = 32'h00312413; // XORI  x8, x2, 3       ; x8 = x2 ^ 3 = 8 ^ 3 = 11
        mem[5] = 32'h00113613; // ORI   x12, x2, 1      ; x12 = x2 | 1 = 9
        mem[6] = 32'h00114613; // ANDI  x12, x2, 1      ; x12 = x2 & 1 = 0
        mem[7] = 32'h00115513; // SLLI  x10, x2, 1      ; x10 = x2 << 1 = 16
        mem[8] = 32'h00116513; // SRLI  x10, x2, 1      ; x10 = x2 >> 1 = 4
        mem[9] = 32'h40117513; // SRAI  x10, x2, 1      ; x10 = arithmetic right shift x2 >> 1 = 4

//    mem[0] = 32'h00500093; // ADDI x1, x0, 5
//    mem[1] = 32'h00500113; // ADDI x2, x0, 5
//    mem[2] = 32'h00808263; // BEQ x1, x2, +8  → jump from PC=8 to PC=16
//    mem[3] = 32'h00000013; // NOP (skipped if branch)
//    mem[4] = 32'h00100193; // ADDI x3, x0, 1
//    mem[5] = 32'h00200213; // ADDI x4, x0, 2
////    Expected PC outputs: 0 → 4 → 8 → 16 → 20 → 24
 
    end 
    
    
assign data_out = mem[addr];
endmodule
